module hazardUnit(input  logic [4:0]  match,
					  input  logic	RegWriteM, RegWriteW, MemtoRegE, 
					  output logic [1:0]  forwardAE, forwardBE,
					  output logic stallD, stallF, flushD, flushE);					 
endmodule 